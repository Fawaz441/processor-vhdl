library ieee;
use ieee.std_logic_1164.all;

entity processor is
    Port(clk: in std_logic;
        value: out std_logic_vector (7 downto 0)
    );

end processor;

architecture Behavioral of processor is

    begin

end Behavioral;